// eth_nios_v2.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module eth_nios_v2 (
		input  wire        clk_clk,                                     //                                   clk.clk
		output wire        eth_tse_0_mac_mdio_connection_mdc,           //         eth_tse_0_mac_mdio_connection.mdc
		input  wire        eth_tse_0_mac_mdio_connection_mdio_in,       //                                      .mdio_in
		output wire        eth_tse_0_mac_mdio_connection_mdio_out,      //                                      .mdio_out
		output wire        eth_tse_0_mac_mdio_connection_mdio_oen,      //                                      .mdio_oen
		output wire        eth_tse_0_mac_misc_connection_magic_wakeup,  //         eth_tse_0_mac_misc_connection.magic_wakeup
		input  wire        eth_tse_0_mac_misc_connection_magic_sleep_n, //                                      .magic_sleep_n
		input  wire        eth_tse_0_mac_misc_connection_ff_tx_crc_fwd, //                                      .ff_tx_crc_fwd
		output wire        eth_tse_0_mac_misc_connection_ff_tx_septy,   //                                      .ff_tx_septy
		output wire        eth_tse_0_mac_misc_connection_tx_ff_uflow,   //                                      .tx_ff_uflow
		output wire        eth_tse_0_mac_misc_connection_ff_tx_a_full,  //                                      .ff_tx_a_full
		output wire        eth_tse_0_mac_misc_connection_ff_tx_a_empty, //                                      .ff_tx_a_empty
		output wire [17:0] eth_tse_0_mac_misc_connection_rx_err_stat,   //                                      .rx_err_stat
		output wire [3:0]  eth_tse_0_mac_misc_connection_rx_frm_type,   //                                      .rx_frm_type
		output wire        eth_tse_0_mac_misc_connection_ff_rx_dsav,    //                                      .ff_rx_dsav
		output wire        eth_tse_0_mac_misc_connection_ff_rx_a_full,  //                                      .ff_rx_a_full
		output wire        eth_tse_0_mac_misc_connection_ff_rx_a_empty, //                                      .ff_rx_a_empty
		input  wire [3:0]  eth_tse_0_mac_rgmii_connection_rgmii_in,     //        eth_tse_0_mac_rgmii_connection.rgmii_in
		output wire [3:0]  eth_tse_0_mac_rgmii_connection_rgmii_out,    //                                      .rgmii_out
		input  wire        eth_tse_0_mac_rgmii_connection_rx_control,   //                                      .rx_control
		output wire        eth_tse_0_mac_rgmii_connection_tx_control,   //                                      .tx_control
		input  wire        eth_tse_0_mac_status_connection_set_10,      //       eth_tse_0_mac_status_connection.set_10
		input  wire        eth_tse_0_mac_status_connection_set_1000,    //                                      .set_1000
		output wire        eth_tse_0_mac_status_connection_eth_mode,    //                                      .eth_mode
		output wire        eth_tse_0_mac_status_connection_ena_10,      //                                      .ena_10
		input  wire        eth_tse_0_pcs_mac_rx_clock_connection_clk,   // eth_tse_0_pcs_mac_rx_clock_connection.clk
		input  wire        eth_tse_0_pcs_mac_tx_clock_connection_clk,   // eth_tse_0_pcs_mac_tx_clock_connection.clk
		input  wire        irq_eth_input_export,                        //                         irq_eth_input.export
		input  wire        rx_tx_buf_clk2_clk,                          //                        rx_tx_buf_clk2.clk
		input  wire        rx_tx_buf_reset2_reset,                      //                      rx_tx_buf_reset2.reset
		input  wire        rx_tx_buf_reset2_reset_req,                  //                                      .reset_req
		input  wire [10:0] rx_tx_buf_s2_address,                        //                          rx_tx_buf_s2.address
		input  wire        rx_tx_buf_s2_chipselect,                     //                                      .chipselect
		input  wire        rx_tx_buf_s2_clken,                          //                                      .clken
		input  wire        rx_tx_buf_s2_write,                          //                                      .write
		output wire [7:0]  rx_tx_buf_s2_readdata,                       //                                      .readdata
		input  wire [7:0]  rx_tx_buf_s2_writedata                       //                                      .writedata
	);

	wire         tx_dma_out_valid;                                            // tx_dma:out_valid -> tse:ff_tx_wren
	wire   [7:0] tx_dma_out_data;                                             // tx_dma:out_data -> tse:ff_tx_data
	wire         tx_dma_out_ready;                                            // tse:ff_tx_rdy -> tx_dma:out_ready
	wire         tx_dma_out_startofpacket;                                    // tx_dma:out_startofpacket -> tse:ff_tx_sop
	wire         tx_dma_out_endofpacket;                                      // tx_dma:out_endofpacket -> tse:ff_tx_eop
	wire         tx_dma_out_error;                                            // tx_dma:out_error -> tse:ff_tx_err
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in0, rst_controller:reset_in1]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [14:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire         rx_dma_m_write_waitrequest;                                  // mm_interconnect_0:rx_dma_m_write_waitrequest -> rx_dma:m_write_waitrequest
	wire  [31:0] rx_dma_m_write_address;                                      // rx_dma:m_write_address -> mm_interconnect_0:rx_dma_m_write_address
	wire         rx_dma_m_write_write;                                        // rx_dma:m_write_write -> mm_interconnect_0:rx_dma_m_write_write
	wire   [7:0] rx_dma_m_write_writedata;                                    // rx_dma:m_write_writedata -> mm_interconnect_0:rx_dma_m_write_writedata
	wire   [7:0] tx_dma_m_read_readdata;                                      // mm_interconnect_0:tx_dma_m_read_readdata -> tx_dma:m_read_readdata
	wire         tx_dma_m_read_waitrequest;                                   // mm_interconnect_0:tx_dma_m_read_waitrequest -> tx_dma:m_read_waitrequest
	wire  [31:0] tx_dma_m_read_address;                                       // tx_dma:m_read_address -> mm_interconnect_0:tx_dma_m_read_address
	wire         tx_dma_m_read_read;                                          // tx_dma:m_read_read -> mm_interconnect_0:tx_dma_m_read_read
	wire         tx_dma_m_read_readdatavalid;                                 // mm_interconnect_0:tx_dma_m_read_readdatavalid -> tx_dma:m_read_readdatavalid
	wire  [31:0] rx_dma_descriptor_read_readdata;                             // mm_interconnect_0:rx_dma_descriptor_read_readdata -> rx_dma:descriptor_read_readdata
	wire         rx_dma_descriptor_read_waitrequest;                          // mm_interconnect_0:rx_dma_descriptor_read_waitrequest -> rx_dma:descriptor_read_waitrequest
	wire  [31:0] rx_dma_descriptor_read_address;                              // rx_dma:descriptor_read_address -> mm_interconnect_0:rx_dma_descriptor_read_address
	wire         rx_dma_descriptor_read_read;                                 // rx_dma:descriptor_read_read -> mm_interconnect_0:rx_dma_descriptor_read_read
	wire         rx_dma_descriptor_read_readdatavalid;                        // mm_interconnect_0:rx_dma_descriptor_read_readdatavalid -> rx_dma:descriptor_read_readdatavalid
	wire  [31:0] tx_dma_descriptor_read_readdata;                             // mm_interconnect_0:tx_dma_descriptor_read_readdata -> tx_dma:descriptor_read_readdata
	wire         tx_dma_descriptor_read_waitrequest;                          // mm_interconnect_0:tx_dma_descriptor_read_waitrequest -> tx_dma:descriptor_read_waitrequest
	wire  [31:0] tx_dma_descriptor_read_address;                              // tx_dma:descriptor_read_address -> mm_interconnect_0:tx_dma_descriptor_read_address
	wire         tx_dma_descriptor_read_read;                                 // tx_dma:descriptor_read_read -> mm_interconnect_0:tx_dma_descriptor_read_read
	wire         tx_dma_descriptor_read_readdatavalid;                        // mm_interconnect_0:tx_dma_descriptor_read_readdatavalid -> tx_dma:descriptor_read_readdatavalid
	wire         rx_dma_descriptor_write_waitrequest;                         // mm_interconnect_0:rx_dma_descriptor_write_waitrequest -> rx_dma:descriptor_write_waitrequest
	wire  [31:0] rx_dma_descriptor_write_address;                             // rx_dma:descriptor_write_address -> mm_interconnect_0:rx_dma_descriptor_write_address
	wire         rx_dma_descriptor_write_write;                               // rx_dma:descriptor_write_write -> mm_interconnect_0:rx_dma_descriptor_write_write
	wire  [31:0] rx_dma_descriptor_write_writedata;                           // rx_dma:descriptor_write_writedata -> mm_interconnect_0:rx_dma_descriptor_write_writedata
	wire         tx_dma_descriptor_write_waitrequest;                         // mm_interconnect_0:tx_dma_descriptor_write_waitrequest -> tx_dma:descriptor_write_waitrequest
	wire  [31:0] tx_dma_descriptor_write_address;                             // tx_dma:descriptor_write_address -> mm_interconnect_0:tx_dma_descriptor_write_address
	wire         tx_dma_descriptor_write_write;                               // tx_dma:descriptor_write_write -> mm_interconnect_0:tx_dma_descriptor_write_write
	wire  [31:0] tx_dma_descriptor_write_writedata;                           // tx_dma:descriptor_write_writedata -> mm_interconnect_0:tx_dma_descriptor_write_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [14:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_tse_control_port_readdata;                 // tse:reg_data_out -> mm_interconnect_0:tse_control_port_readdata
	wire         mm_interconnect_0_tse_control_port_waitrequest;              // tse:reg_busy -> mm_interconnect_0:tse_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_control_port_address;                  // mm_interconnect_0:tse_control_port_address -> tse:reg_addr
	wire         mm_interconnect_0_tse_control_port_read;                     // mm_interconnect_0:tse_control_port_read -> tse:reg_rd
	wire         mm_interconnect_0_tse_control_port_write;                    // mm_interconnect_0:tse_control_port_write -> tse:reg_wr
	wire  [31:0] mm_interconnect_0_tse_control_port_writedata;                // mm_interconnect_0:tse_control_port_writedata -> tse:reg_data_in
	wire         mm_interconnect_0_tx_dma_csr_chipselect;                     // mm_interconnect_0:tx_dma_csr_chipselect -> tx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_tx_dma_csr_readdata;                       // tx_dma:csr_readdata -> mm_interconnect_0:tx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_tx_dma_csr_address;                        // mm_interconnect_0:tx_dma_csr_address -> tx_dma:csr_address
	wire         mm_interconnect_0_tx_dma_csr_read;                           // mm_interconnect_0:tx_dma_csr_read -> tx_dma:csr_read
	wire         mm_interconnect_0_tx_dma_csr_write;                          // mm_interconnect_0:tx_dma_csr_write -> tx_dma:csr_write
	wire  [31:0] mm_interconnect_0_tx_dma_csr_writedata;                      // mm_interconnect_0:tx_dma_csr_writedata -> tx_dma:csr_writedata
	wire         mm_interconnect_0_rx_dma_csr_chipselect;                     // mm_interconnect_0:rx_dma_csr_chipselect -> rx_dma:csr_chipselect
	wire  [31:0] mm_interconnect_0_rx_dma_csr_readdata;                       // rx_dma:csr_readdata -> mm_interconnect_0:rx_dma_csr_readdata
	wire   [3:0] mm_interconnect_0_rx_dma_csr_address;                        // mm_interconnect_0:rx_dma_csr_address -> rx_dma:csr_address
	wire         mm_interconnect_0_rx_dma_csr_read;                           // mm_interconnect_0:rx_dma_csr_read -> rx_dma:csr_read
	wire         mm_interconnect_0_rx_dma_csr_write;                          // mm_interconnect_0:rx_dma_csr_write -> rx_dma:csr_write
	wire  [31:0] mm_interconnect_0_rx_dma_csr_writedata;                      // mm_interconnect_0:rx_dma_csr_writedata -> rx_dma:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_system_ram_s1_chipselect;                  // mm_interconnect_0:system_ram_s1_chipselect -> system_ram:chipselect
	wire  [31:0] mm_interconnect_0_system_ram_s1_readdata;                    // system_ram:readdata -> mm_interconnect_0:system_ram_s1_readdata
	wire  [10:0] mm_interconnect_0_system_ram_s1_address;                     // mm_interconnect_0:system_ram_s1_address -> system_ram:address
	wire   [3:0] mm_interconnect_0_system_ram_s1_byteenable;                  // mm_interconnect_0:system_ram_s1_byteenable -> system_ram:byteenable
	wire         mm_interconnect_0_system_ram_s1_write;                       // mm_interconnect_0:system_ram_s1_write -> system_ram:write
	wire  [31:0] mm_interconnect_0_system_ram_s1_writedata;                   // mm_interconnect_0:system_ram_s1_writedata -> system_ram:writedata
	wire         mm_interconnect_0_system_ram_s1_clken;                       // mm_interconnect_0:system_ram_s1_clken -> system_ram:clken
	wire         mm_interconnect_0_header_ram_s1_chipselect;                  // mm_interconnect_0:header_ram_s1_chipselect -> header_ram:chipselect
	wire   [7:0] mm_interconnect_0_header_ram_s1_readdata;                    // header_ram:readdata -> mm_interconnect_0:header_ram_s1_readdata
	wire   [7:0] mm_interconnect_0_header_ram_s1_address;                     // mm_interconnect_0:header_ram_s1_address -> header_ram:address
	wire         mm_interconnect_0_header_ram_s1_write;                       // mm_interconnect_0:header_ram_s1_write -> header_ram:write
	wire   [7:0] mm_interconnect_0_header_ram_s1_writedata;                   // mm_interconnect_0:header_ram_s1_writedata -> header_ram:writedata
	wire         mm_interconnect_0_header_ram_s1_clken;                       // mm_interconnect_0:header_ram_s1_clken -> header_ram:clken
	wire         mm_interconnect_0_timer_0_s1_chipselect;                     // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                       // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                        // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                          // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                      // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_rx_buf_ram_s1_chipselect;                  // mm_interconnect_0:rx_buf_ram_s1_chipselect -> rx_buf_ram:chipselect
	wire   [7:0] mm_interconnect_0_rx_buf_ram_s1_readdata;                    // rx_buf_ram:readdata -> mm_interconnect_0:rx_buf_ram_s1_readdata
	wire   [8:0] mm_interconnect_0_rx_buf_ram_s1_address;                     // mm_interconnect_0:rx_buf_ram_s1_address -> rx_buf_ram:address
	wire         mm_interconnect_0_rx_buf_ram_s1_write;                       // mm_interconnect_0:rx_buf_ram_s1_write -> rx_buf_ram:write
	wire   [7:0] mm_interconnect_0_rx_buf_ram_s1_writedata;                   // mm_interconnect_0:rx_buf_ram_s1_writedata -> rx_buf_ram:writedata
	wire         mm_interconnect_0_rx_buf_ram_s1_clken;                       // mm_interconnect_0:rx_buf_ram_s1_clken -> rx_buf_ram:clken
	wire         mm_interconnect_0_eth_irq_pio_s1_chipselect;                 // mm_interconnect_0:eth_irq_pio_s1_chipselect -> eth_irq_pio:chipselect
	wire  [31:0] mm_interconnect_0_eth_irq_pio_s1_readdata;                   // eth_irq_pio:readdata -> mm_interconnect_0:eth_irq_pio_s1_readdata
	wire   [1:0] mm_interconnect_0_eth_irq_pio_s1_address;                    // mm_interconnect_0:eth_irq_pio_s1_address -> eth_irq_pio:address
	wire         mm_interconnect_0_eth_irq_pio_s1_write;                      // mm_interconnect_0:eth_irq_pio_s1_write -> eth_irq_pio:write_n
	wire  [31:0] mm_interconnect_0_eth_irq_pio_s1_writedata;                  // mm_interconnect_0:eth_irq_pio_s1_writedata -> eth_irq_pio:writedata
	wire         mm_interconnect_0_tx_buff_ram_s1_chipselect;                 // mm_interconnect_0:tx_buff_ram_s1_chipselect -> tx_buff_ram:chipselect
	wire   [7:0] mm_interconnect_0_tx_buff_ram_s1_readdata;                   // tx_buff_ram:readdata -> mm_interconnect_0:tx_buff_ram_s1_readdata
	wire  [10:0] mm_interconnect_0_tx_buff_ram_s1_address;                    // mm_interconnect_0:tx_buff_ram_s1_address -> tx_buff_ram:address
	wire         mm_interconnect_0_tx_buff_ram_s1_write;                      // mm_interconnect_0:tx_buff_ram_s1_write -> tx_buff_ram:write
	wire   [7:0] mm_interconnect_0_tx_buff_ram_s1_writedata;                  // mm_interconnect_0:tx_buff_ram_s1_writedata -> tx_buff_ram:writedata
	wire         mm_interconnect_0_tx_buff_ram_s1_clken;                      // mm_interconnect_0:tx_buff_ram_s1_clken -> tx_buff_ram:clken
	wire         irq_mapper_receiver0_irq;                                    // rx_dma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                    // tx_dma:csr_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                    // timer_0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                    // eth_irq_pio:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         tse_receive_valid;                                           // tse:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire   [7:0] tse_receive_data;                                            // tse:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_receive_ready;                                           // avalon_st_adapter:in_0_ready -> tse:ff_rx_rdy
	wire         tse_receive_startofpacket;                                   // tse:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_receive_endofpacket;                                     // tse:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_receive_error;                                           // tse:rx_err -> avalon_st_adapter:in_0_error
	wire         avalon_st_adapter_out_0_valid;                               // avalon_st_adapter:out_0_valid -> rx_dma:in_valid
	wire   [7:0] avalon_st_adapter_out_0_data;                                // avalon_st_adapter:out_0_data -> rx_dma:in_data
	wire         avalon_st_adapter_out_0_ready;                               // rx_dma:in_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                       // avalon_st_adapter:out_0_startofpacket -> rx_dma:in_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                         // avalon_st_adapter:out_0_endofpacket -> rx_dma:in_endofpacket
	wire         avalon_st_adapter_out_0_error;                               // avalon_st_adapter:out_0_error -> rx_dma:in_error
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, eth_irq_pio:reset_n, header_ram:reset, irq_mapper:reset, jtag_uart_0:rst_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, rst_translator:in_reset, rx_buf_ram:reset, rx_dma:system_reset_n, system_ram:reset, timer_0:reset_n, tse:reset, tx_buff_ram:reset, tx_dma:system_reset_n]
	wire         rst_controller_reset_out_reset_req;                          // rst_controller:reset_req -> [header_ram:reset_req, nios2_gen2_0:reset_req, rst_translator:reset_req_in, rx_buf_ram:reset_req, system_ram:reset_req, tx_buff_ram:reset_req]

	eth_nios_v2_eth_irq_pio eth_irq_pio (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_eth_irq_pio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_eth_irq_pio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_eth_irq_pio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_eth_irq_pio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_eth_irq_pio_s1_readdata),   //                    .readdata
		.in_port    (irq_eth_input_export),                        // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                     //                 irq.irq
	);

	eth_nios_v2_header_ram header_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_header_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_header_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_header_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_header_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_header_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_header_ram_s1_writedata),  //       .writedata
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	eth_nios_v2_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                                     //               irq.irq
	);

	eth_nios_v2_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	eth_nios_v2_rx_buf_ram rx_buf_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_rx_buf_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_rx_buf_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_rx_buf_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_rx_buf_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_rx_buf_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_rx_buf_ram_s1_writedata),  //       .writedata
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	eth_nios_v2_rx_dma rx_dma (
		.clk                           (clk_clk),                                 //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),         //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_rx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_rx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_rx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_rx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_rx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_rx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (rx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (rx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (rx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (rx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (rx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (rx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (rx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (rx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (rx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                //          csr_irq.irq
		.in_startofpacket              (avalon_st_adapter_out_0_startofpacket),   //               in.startofpacket
		.in_endofpacket                (avalon_st_adapter_out_0_endofpacket),     //                 .endofpacket
		.in_data                       (avalon_st_adapter_out_0_data),            //                 .data
		.in_valid                      (avalon_st_adapter_out_0_valid),           //                 .valid
		.in_ready                      (avalon_st_adapter_out_0_ready),           //                 .ready
		.in_error                      (avalon_st_adapter_out_0_error),           //                 .error
		.m_write_waitrequest           (rx_dma_m_write_waitrequest),              //          m_write.waitrequest
		.m_write_address               (rx_dma_m_write_address),                  //                 .address
		.m_write_write                 (rx_dma_m_write_write),                    //                 .write
		.m_write_writedata             (rx_dma_m_write_writedata)                 //                 .writedata
	);

	eth_nios_v2_system_ram system_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_system_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_system_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_system_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_system_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_system_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_system_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_system_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),         //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	eth_nios_v2_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	eth_nios_v2_tse tse (
		.clk           (clk_clk),                                        // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                 //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (eth_tse_0_pcs_mac_tx_clock_connection_clk),      //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (eth_tse_0_pcs_mac_rx_clock_connection_clk),      //   pcs_mac_rx_clock_connection.clk
		.set_10        (eth_tse_0_mac_status_connection_set_10),         //         mac_status_connection.set_10
		.set_1000      (eth_tse_0_mac_status_connection_set_1000),       //                              .set_1000
		.eth_mode      (eth_tse_0_mac_status_connection_eth_mode),       //                              .eth_mode
		.ena_10        (eth_tse_0_mac_status_connection_ena_10),         //                              .ena_10
		.rgmii_in      (eth_tse_0_mac_rgmii_connection_rgmii_in),        //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (eth_tse_0_mac_rgmii_connection_rgmii_out),       //                              .rgmii_out
		.rx_control    (eth_tse_0_mac_rgmii_connection_rx_control),      //                              .rx_control
		.tx_control    (eth_tse_0_mac_rgmii_connection_tx_control),      //                              .tx_control
		.ff_rx_clk     (clk_clk),                                        //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                        //     transmit_clock_connection.clk
		.ff_rx_data    (tse_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_receive_error),                              //                              .error
		.ff_rx_rdy     (tse_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_receive_valid),                              //                              .valid
		.ff_tx_data    (tx_dma_out_data),                                //                      transmit.data
		.ff_tx_eop     (tx_dma_out_endofpacket),                         //                              .endofpacket
		.ff_tx_err     (tx_dma_out_error),                               //                              .error
		.ff_tx_rdy     (tx_dma_out_ready),                               //                              .ready
		.ff_tx_sop     (tx_dma_out_startofpacket),                       //                              .startofpacket
		.ff_tx_wren    (tx_dma_out_valid),                               //                              .valid
		.mdc           (eth_tse_0_mac_mdio_connection_mdc),              //           mac_mdio_connection.mdc
		.mdio_in       (eth_tse_0_mac_mdio_connection_mdio_in),          //                              .mdio_in
		.mdio_out      (eth_tse_0_mac_mdio_connection_mdio_out),         //                              .mdio_out
		.mdio_oen      (eth_tse_0_mac_mdio_connection_mdio_oen),         //                              .mdio_oen
		.magic_wakeup  (eth_tse_0_mac_misc_connection_magic_wakeup),     //           mac_misc_connection.magic_wakeup
		.magic_sleep_n (eth_tse_0_mac_misc_connection_magic_sleep_n),    //                              .magic_sleep_n
		.ff_tx_crc_fwd (eth_tse_0_mac_misc_connection_ff_tx_crc_fwd),    //                              .ff_tx_crc_fwd
		.ff_tx_septy   (eth_tse_0_mac_misc_connection_ff_tx_septy),      //                              .ff_tx_septy
		.tx_ff_uflow   (eth_tse_0_mac_misc_connection_tx_ff_uflow),      //                              .tx_ff_uflow
		.ff_tx_a_full  (eth_tse_0_mac_misc_connection_ff_tx_a_full),     //                              .ff_tx_a_full
		.ff_tx_a_empty (eth_tse_0_mac_misc_connection_ff_tx_a_empty),    //                              .ff_tx_a_empty
		.rx_err_stat   (eth_tse_0_mac_misc_connection_rx_err_stat),      //                              .rx_err_stat
		.rx_frm_type   (eth_tse_0_mac_misc_connection_rx_frm_type),      //                              .rx_frm_type
		.ff_rx_dsav    (eth_tse_0_mac_misc_connection_ff_rx_dsav),       //                              .ff_rx_dsav
		.ff_rx_a_full  (eth_tse_0_mac_misc_connection_ff_rx_a_full),     //                              .ff_rx_a_full
		.ff_rx_a_empty (eth_tse_0_mac_misc_connection_ff_rx_a_empty)     //                              .ff_rx_a_empty
	);

	eth_nios_v2_tx_buff_ram tx_buff_ram (
		.clk         (clk_clk),                                     //   clk1.clk
		.address     (mm_interconnect_0_tx_buff_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_tx_buff_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_tx_buff_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_tx_buff_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_tx_buff_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_tx_buff_ram_s1_writedata),  //       .writedata
		.reset       (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),          //       .reset_req
		.address2    (rx_tx_buf_s2_address),                        //     s2.address
		.chipselect2 (rx_tx_buf_s2_chipselect),                     //       .chipselect
		.clken2      (rx_tx_buf_s2_clken),                          //       .clken
		.write2      (rx_tx_buf_s2_write),                          //       .write
		.readdata2   (rx_tx_buf_s2_readdata),                       //       .readdata
		.writedata2  (rx_tx_buf_s2_writedata),                      //       .writedata
		.clk2        (rx_tx_buf_clk2_clk),                          //   clk2.clk
		.reset2      (rx_tx_buf_reset2_reset),                      // reset2.reset
		.reset_req2  (rx_tx_buf_reset2_reset_req),                  //       .reset_req
		.freeze      (1'b0)                                         // (terminated)
	);

	eth_nios_v2_tx_dma tx_dma (
		.clk                           (clk_clk),                                 //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),         //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_tx_dma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_tx_dma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_tx_dma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_tx_dma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_tx_dma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_tx_dma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (tx_dma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (tx_dma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (tx_dma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (tx_dma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (tx_dma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (tx_dma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (tx_dma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (tx_dma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (tx_dma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver1_irq),                //          csr_irq.irq
		.m_read_readdata               (tx_dma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (tx_dma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (tx_dma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (tx_dma_m_read_address),                   //                 .address
		.m_read_read                   (tx_dma_m_read_read),                      //                 .read
		.out_data                      (tx_dma_out_data),                         //              out.data
		.out_valid                     (tx_dma_out_valid),                        //                 .valid
		.out_ready                     (tx_dma_out_ready),                        //                 .ready
		.out_endofpacket               (tx_dma_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (tx_dma_out_startofpacket),                //                 .startofpacket
		.out_error                     (tx_dma_out_error)                         //                 .error
	);

	eth_nios_v2_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                              // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_readdatavalid         (nios2_gen2_0_data_master_readdatavalid),                      //                                         .readdatavalid
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.nios2_gen2_0_instruction_master_readdatavalid  (nios2_gen2_0_instruction_master_readdatavalid),               //                                         .readdatavalid
		.rx_dma_descriptor_read_address                 (rx_dma_descriptor_read_address),                              //                   rx_dma_descriptor_read.address
		.rx_dma_descriptor_read_waitrequest             (rx_dma_descriptor_read_waitrequest),                          //                                         .waitrequest
		.rx_dma_descriptor_read_read                    (rx_dma_descriptor_read_read),                                 //                                         .read
		.rx_dma_descriptor_read_readdata                (rx_dma_descriptor_read_readdata),                             //                                         .readdata
		.rx_dma_descriptor_read_readdatavalid           (rx_dma_descriptor_read_readdatavalid),                        //                                         .readdatavalid
		.rx_dma_descriptor_write_address                (rx_dma_descriptor_write_address),                             //                  rx_dma_descriptor_write.address
		.rx_dma_descriptor_write_waitrequest            (rx_dma_descriptor_write_waitrequest),                         //                                         .waitrequest
		.rx_dma_descriptor_write_write                  (rx_dma_descriptor_write_write),                               //                                         .write
		.rx_dma_descriptor_write_writedata              (rx_dma_descriptor_write_writedata),                           //                                         .writedata
		.rx_dma_m_write_address                         (rx_dma_m_write_address),                                      //                           rx_dma_m_write.address
		.rx_dma_m_write_waitrequest                     (rx_dma_m_write_waitrequest),                                  //                                         .waitrequest
		.rx_dma_m_write_write                           (rx_dma_m_write_write),                                        //                                         .write
		.rx_dma_m_write_writedata                       (rx_dma_m_write_writedata),                                    //                                         .writedata
		.tx_dma_descriptor_read_address                 (tx_dma_descriptor_read_address),                              //                   tx_dma_descriptor_read.address
		.tx_dma_descriptor_read_waitrequest             (tx_dma_descriptor_read_waitrequest),                          //                                         .waitrequest
		.tx_dma_descriptor_read_read                    (tx_dma_descriptor_read_read),                                 //                                         .read
		.tx_dma_descriptor_read_readdata                (tx_dma_descriptor_read_readdata),                             //                                         .readdata
		.tx_dma_descriptor_read_readdatavalid           (tx_dma_descriptor_read_readdatavalid),                        //                                         .readdatavalid
		.tx_dma_descriptor_write_address                (tx_dma_descriptor_write_address),                             //                  tx_dma_descriptor_write.address
		.tx_dma_descriptor_write_waitrequest            (tx_dma_descriptor_write_waitrequest),                         //                                         .waitrequest
		.tx_dma_descriptor_write_write                  (tx_dma_descriptor_write_write),                               //                                         .write
		.tx_dma_descriptor_write_writedata              (tx_dma_descriptor_write_writedata),                           //                                         .writedata
		.tx_dma_m_read_address                          (tx_dma_m_read_address),                                       //                            tx_dma_m_read.address
		.tx_dma_m_read_waitrequest                      (tx_dma_m_read_waitrequest),                                   //                                         .waitrequest
		.tx_dma_m_read_read                             (tx_dma_m_read_read),                                          //                                         .read
		.tx_dma_m_read_readdata                         (tx_dma_m_read_readdata),                                      //                                         .readdata
		.tx_dma_m_read_readdatavalid                    (tx_dma_m_read_readdatavalid),                                 //                                         .readdatavalid
		.eth_irq_pio_s1_address                         (mm_interconnect_0_eth_irq_pio_s1_address),                    //                           eth_irq_pio_s1.address
		.eth_irq_pio_s1_write                           (mm_interconnect_0_eth_irq_pio_s1_write),                      //                                         .write
		.eth_irq_pio_s1_readdata                        (mm_interconnect_0_eth_irq_pio_s1_readdata),                   //                                         .readdata
		.eth_irq_pio_s1_writedata                       (mm_interconnect_0_eth_irq_pio_s1_writedata),                  //                                         .writedata
		.eth_irq_pio_s1_chipselect                      (mm_interconnect_0_eth_irq_pio_s1_chipselect),                 //                                         .chipselect
		.header_ram_s1_address                          (mm_interconnect_0_header_ram_s1_address),                     //                            header_ram_s1.address
		.header_ram_s1_write                            (mm_interconnect_0_header_ram_s1_write),                       //                                         .write
		.header_ram_s1_readdata                         (mm_interconnect_0_header_ram_s1_readdata),                    //                                         .readdata
		.header_ram_s1_writedata                        (mm_interconnect_0_header_ram_s1_writedata),                   //                                         .writedata
		.header_ram_s1_chipselect                       (mm_interconnect_0_header_ram_s1_chipselect),                  //                                         .chipselect
		.header_ram_s1_clken                            (mm_interconnect_0_header_ram_s1_clken),                       //                                         .clken
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.rx_buf_ram_s1_address                          (mm_interconnect_0_rx_buf_ram_s1_address),                     //                            rx_buf_ram_s1.address
		.rx_buf_ram_s1_write                            (mm_interconnect_0_rx_buf_ram_s1_write),                       //                                         .write
		.rx_buf_ram_s1_readdata                         (mm_interconnect_0_rx_buf_ram_s1_readdata),                    //                                         .readdata
		.rx_buf_ram_s1_writedata                        (mm_interconnect_0_rx_buf_ram_s1_writedata),                   //                                         .writedata
		.rx_buf_ram_s1_chipselect                       (mm_interconnect_0_rx_buf_ram_s1_chipselect),                  //                                         .chipselect
		.rx_buf_ram_s1_clken                            (mm_interconnect_0_rx_buf_ram_s1_clken),                       //                                         .clken
		.rx_dma_csr_address                             (mm_interconnect_0_rx_dma_csr_address),                        //                               rx_dma_csr.address
		.rx_dma_csr_write                               (mm_interconnect_0_rx_dma_csr_write),                          //                                         .write
		.rx_dma_csr_read                                (mm_interconnect_0_rx_dma_csr_read),                           //                                         .read
		.rx_dma_csr_readdata                            (mm_interconnect_0_rx_dma_csr_readdata),                       //                                         .readdata
		.rx_dma_csr_writedata                           (mm_interconnect_0_rx_dma_csr_writedata),                      //                                         .writedata
		.rx_dma_csr_chipselect                          (mm_interconnect_0_rx_dma_csr_chipselect),                     //                                         .chipselect
		.system_ram_s1_address                          (mm_interconnect_0_system_ram_s1_address),                     //                            system_ram_s1.address
		.system_ram_s1_write                            (mm_interconnect_0_system_ram_s1_write),                       //                                         .write
		.system_ram_s1_readdata                         (mm_interconnect_0_system_ram_s1_readdata),                    //                                         .readdata
		.system_ram_s1_writedata                        (mm_interconnect_0_system_ram_s1_writedata),                   //                                         .writedata
		.system_ram_s1_byteenable                       (mm_interconnect_0_system_ram_s1_byteenable),                  //                                         .byteenable
		.system_ram_s1_chipselect                       (mm_interconnect_0_system_ram_s1_chipselect),                  //                                         .chipselect
		.system_ram_s1_clken                            (mm_interconnect_0_system_ram_s1_clken),                       //                                         .clken
		.timer_0_s1_address                             (mm_interconnect_0_timer_0_s1_address),                        //                               timer_0_s1.address
		.timer_0_s1_write                               (mm_interconnect_0_timer_0_s1_write),                          //                                         .write
		.timer_0_s1_readdata                            (mm_interconnect_0_timer_0_s1_readdata),                       //                                         .readdata
		.timer_0_s1_writedata                           (mm_interconnect_0_timer_0_s1_writedata),                      //                                         .writedata
		.timer_0_s1_chipselect                          (mm_interconnect_0_timer_0_s1_chipselect),                     //                                         .chipselect
		.tse_control_port_address                       (mm_interconnect_0_tse_control_port_address),                  //                         tse_control_port.address
		.tse_control_port_write                         (mm_interconnect_0_tse_control_port_write),                    //                                         .write
		.tse_control_port_read                          (mm_interconnect_0_tse_control_port_read),                     //                                         .read
		.tse_control_port_readdata                      (mm_interconnect_0_tse_control_port_readdata),                 //                                         .readdata
		.tse_control_port_writedata                     (mm_interconnect_0_tse_control_port_writedata),                //                                         .writedata
		.tse_control_port_waitrequest                   (mm_interconnect_0_tse_control_port_waitrequest),              //                                         .waitrequest
		.tx_buff_ram_s1_address                         (mm_interconnect_0_tx_buff_ram_s1_address),                    //                           tx_buff_ram_s1.address
		.tx_buff_ram_s1_write                           (mm_interconnect_0_tx_buff_ram_s1_write),                      //                                         .write
		.tx_buff_ram_s1_readdata                        (mm_interconnect_0_tx_buff_ram_s1_readdata),                   //                                         .readdata
		.tx_buff_ram_s1_writedata                       (mm_interconnect_0_tx_buff_ram_s1_writedata),                  //                                         .writedata
		.tx_buff_ram_s1_chipselect                      (mm_interconnect_0_tx_buff_ram_s1_chipselect),                 //                                         .chipselect
		.tx_buff_ram_s1_clken                           (mm_interconnect_0_tx_buff_ram_s1_clken),                      //                                         .clken
		.tx_dma_csr_address                             (mm_interconnect_0_tx_dma_csr_address),                        //                               tx_dma_csr.address
		.tx_dma_csr_write                               (mm_interconnect_0_tx_dma_csr_write),                          //                                         .write
		.tx_dma_csr_read                                (mm_interconnect_0_tx_dma_csr_read),                           //                                         .read
		.tx_dma_csr_readdata                            (mm_interconnect_0_tx_dma_csr_readdata),                       //                                         .readdata
		.tx_dma_csr_writedata                           (mm_interconnect_0_tx_dma_csr_writedata),                      //                                         .writedata
		.tx_dma_csr_chipselect                          (mm_interconnect_0_tx_dma_csr_chipselect)                      //                                         .chipselect
	);

	eth_nios_v2_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	eth_nios_v2_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (8),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (8),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (tse_receive_data),                      //     in_0.data
		.in_0_valid          (tse_receive_valid),                     //         .valid
		.in_0_ready          (tse_receive_ready),                     //         .ready
		.in_0_startofpacket  (tse_receive_startofpacket),             //         .startofpacket
		.in_0_endofpacket    (tse_receive_endofpacket),               //         .endofpacket
		.in_0_error          (tse_receive_error),                     //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_0_debug_reset_request_reset), // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
