module DMAcontroller
();



/*                                                                                                                                                                                                                                                                                                                                
	Модули обращаются к DMA контроллеру с запросом на доступ к памяти. Задача контроллера арббитраж запросов.
Арбитраж может проводиться в зависимости от приоритетов, например от чтения с самым высоким приоритетом к записии с 
самым низким приоритетом, от больших транзакций к малым, то есть, приоритет отдается модулю который хочет прочитать большой
объем данных, т.к. чтение позволит системе продолжит совю работу в отличаи от записи.
	Так же возможен арбитраж по времени ожидания, т.е. каждый раз, когда модуль обращается к контроллеру, тот обнуляет счетчик
времени ожидания, приоритет отдается модулю с наибольшим временем ожидания.


	В тот момент, когда контроллер выдает разрешение модулю на обращение к памяти, тот начинает слушать общую шинну данных и шину адреса
либо же контроллер начинает забирать данные из внутренней RAM памяти
	
*/


endmodule
